
module MEM;  
endmodule  

module SC;  
endmodule  

module Xbar;  
endmodule  


module IS;  
    MEM mem1();  
    SC sc1();  
    Xbar xbar1();  
endmodule  


module Top;  
    IS is1();  
endmodule  
